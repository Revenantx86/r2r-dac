module b2t #()();




endmodule